----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    15:51:06 07/24/2016 
-- Design Name: 
-- Module Name:    CONTROL_MEMORY_256x28 - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity CONTROL_MEMORY_256x28 is
Port ( 
	MW : out std_logic;
	MM : out std_logic;
	RW : out std_logic;
	MD : out std_logic;
	FUNC_SEL : out std_logic_vector(4 downto 0);
	MB : out std_logic;
	TB : out std_logic;
	TA : out std_logic;
	TD : out std_logic;
	PL : out std_logic;
	PI : out std_logic;
	IL : out std_logic;
	MC : out std_logic;
	MS_SEL : out std_logic_vector(2 downto 0);
	NA : out std_logic_vector(7 downto 0);
	IN_CAR : in std_logic_vector(7 downto 0));
end CONTROL_MEMORY_256x28;

architecture Behavioral of CONTROL_MEMORY_256x28 is

type mem_array is array(0 to 255) of std_logic_vector(27 downto 0);
begin
	memory_m: process(IN_CAR)
		variable control_mem : mem_array:=(
		------------------------------------------------------------------------------
		------------------------------------------------------------------------------			
		------------------------------------------------------------------------------
		-- INITIALIZE - ADDRESS 0x00 -> 0x03
		------------------------------------------------------------------------------
		------------------------------------------------------------------------------
		------------------------------------------------------------------------------			 
		--NA        MS    MC  IL  PI  PL  TD  TA  TB  MB  FS      MD  RW  MM  MW
		X"01"     &"001"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"10000"&'0'&'0'&'0'&'0', -- 0
		
		X"01"     &"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"10000"&'0'&'0'&'0'&'0', -- 1 
		
		X"02"     &"000"&'0'&'1'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'1'&'0'&'0', -- 2  
		
		X"03"     &"000"&'0'&'0'&'0'&'1'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 3
		------------------------------------------------------------------------------
		------------------------------------------------------------------------------		
		------------------------------------------------------------------------------
		-- END OF INITIALIZE STATE 
		------------------------------------------------------------------------------
		------------------------------------------------------------------------------
		
		------------------------------------------------------------------------------		
		------------------------------------------------------------------------------
		-- GET NEXT INSTRUCTION  -  ADDRESS 0x04 -> 0x06  --
		------------------------------------------------------------------------------
		------------------------------------------------------------------------------
		------------------------------------------------------------------------------
		X"04" 	 &"000"&'0'&'0'&'0'&'0'&'1'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 4		
		X"05"     &"000"&'0'&'0'&'1'&'0'&'1'&'0'&'0'&'0'&"00000"&'0'&'0'&'1'&'0', -- 5  
		X"06"     &"000"&'0'&'1'&'0'&'0'&'1'&'0'&'0'&'0'&"00000"&'0'&'0'&'1'&'0', -- 6 		
		X"07"     &"001"&'1'&'0'&'0'&'0'&'1'&'0'&'0'&'0'&"00000"&'0'&'0'&'1'&'0', -- 7  
		------------------------------------------------------------------------------
		------------------------------------------------------------------------------			
		------------------------------------------------------------------------------
		-- END OF GET NEXT INSTRUCTION 
		------------------------------------------------------------------------------
		------------------------------------------------------------------------------
		
		------------------------------------------------------------------------------		
		------------------------------------------------------------------------------
		-- 
		------------------------------------------------------------------------------
		------------------------------------------------------------------------------
		------------------------------------------------------------------------------		
		X"08"		 &"001"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 8
		X"00"		 &"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 9
		X"00"		 &"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- A 
		------------------------------------------------------------------------------
		------------------------------------------------------------------------------
		------------------------------------------------------------------------------
		-- 
		------------------------------------------------------------------------------
		------------------------------------------------------------------------------
		------------------------------------------------------------------------------		
		X"00"     &"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'1'&'0'&'0'&'0', -- B
		X"00"     &"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'1'&'0'&'0'&'0', -- C    
		X"00"     &"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'1'&'0'&'0'&'0', -- D
		X"00"     &"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'1'&'0'&'0'&'0', -- E     
		X"00"     &"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'1'&'0'&'0'&'0', -- F
	
   	------------------------------------------------------------------
		-- 1					
		------------------------------------------------------------------
		--NA        MS    MC  IL  PI  PL  TD  TA  TB  MB  FS      MD  RW  MM  MW
		X"00" 	 &"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 0		
		X"00"		 &"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 1
		X"00"		 &"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 2
		X"00"		 &"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 3
		
		X"00"		 &"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 4
		X"00"		 &"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 5
		X"00"		 &"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 6
		X"00"		 &"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 7

		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"01000"&'0'&'0'&'0'&'0', -- 8
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"01010"&'0'&'0'&'0'&'0', -- 9
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"01100"&'0'&'0'&'0'&'0', -- A
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"01110"&'0'&'0'&'0'&'0', -- B

		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"10000"&'0'&'0'&'0'&'0', -- C
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"10100"&'0'&'0'&'0'&'0', -- D
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"11000"&'0'&'0'&'0'&'0', -- E
		------------------------------------------------------------------
		-- 1.E				0x1F UNUSED (FOR NOW)
		------------------------------------------------------------------
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- F
		
		------------------------------------------------------------------
		-- 2					YARRR HERE THERE BE AND
		------------------------------------------------------------------
		--NA        MS    MC  IL  PI  PL  TD  TA  TB  MB  FS      MD  RW  MM  MW
		x"20"     &"000"&'0'&'0'&'0'&'0'&'1'&'0'&'0'&'1'&"01000"&'0'&'0'&'0'&'0', -- 0
		x"00"     &"000"&'0'&'0'&'0'&'0'&'1'&'0'&'0'&'1'&"01000"&'0'&'0'&'0'&'0', -- 1
		x"00"		 &"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"01000"&'0'&'1'&'0'&'0', -- 2	
		x"00"		 &"000"&'0'&'0'&'0'&'0'&'1'&'0'&'0'&'0'&"01000"&'0'&'0'&'0'&'0', -- 3
		x"04"		 &"001"&'0'&'0'&'0'&'0'&'1'&'0'&'0'&'0'&"01000"&'0'&'0'&'0'&'0', -- 4
		
		x"25" 	 &"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"01000"&'0'&'0'&'0'&'0', -- 5
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 6
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 7
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 8
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 9
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- A
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- B
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- C
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- D
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- E
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- F
		
		-- ADDRESSES 0x30 -> 0x3F
		--NA        MS    MC  IL  PI  PL  TD  TA  TB  MB  FS      MD  RW  MM  MW
		------------------------------------------------------------------------------		
		------------------------------------------------------------------------------
		-- LDR INSTRUCTION  -  ADDRESS 0x30 -> 0x35
		------------------------------------------------------------------------------
		------------------------------------------------------------------------------
		------------------------------------------------------------------------------
		X"00"		 &"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"11011"&'1'&'0'&'0'&'0', -- 0
		X"00" 	 &"000"&'0'&'0'&'1'&'0'&'0'&'0'&'0'&'0'&"11011"&'1'&'0'&'1'&'0', -- 1		
		X"00"		 &"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"11011"&'1'&'0'&'1'&'0', -- 2
		X"00"		 &"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"11011"&'1'&'1'&'1'&'0', -- 3
		X"00"		 &"000"&'0'&'0'&'0'&'0'&'1'&'0'&'0'&'0'&"11011"&'1'&'0'&'1'&'0', -- 4 
		X"04"		 &"001"&'0'&'0'&'0'&'0'&'1'&'0'&'0'&'0'&"11011"&'1'&'0'&'1'&'0', -- 5 
		------------------------------------------------------------------------------
		------------------------------------------------------------------------------
		------------------------------------------------------------------------------
		-- END OF LDR INSTRUCTION 
		------------------------------------------------------------------------------
		------------------------------------------------------------------------------
		------------------------------------------------------------------------------
		------------------------------------------------------------------------------
		------------------------------------------------------------------------------
		-- STR INSTRUCTION  -  ADDRESS 0x36 -> 0x3D
		------------------------------------------------------------------------------
		------------------------------------------------------------------------------
		X"00"		 &"000"&'0'&'0'&'0'&'0'&'1'&'0'&'0'&'0'&"01111"&'1'&'0'&'1'&'0', -- 6
		X"00"		 &"000"&'0'&'0'&'1'&'0'&'1'&'0'&'0'&'0'&"01111"&'1'&'0'&'1'&'0', -- 7
		X"00"		 &"000"&'0'&'0'&'0'&'0'&'1'&'0'&'0'&'0'&"01111"&'1'&'1'&'1'&'0', -- 8
		X"00"		 &"000"&'0'&'0'&'0'&'0'&'1'&'0'&'0'&'1'&"01111"&'1'&'0'&'1'&'0', -- 9
		X"00"		 &"000"&'0'&'0'&'0'&'0'&'1'&'1'&'0'&'1'&"01111"&'1'&'0'&'0'&'0', -- A
		X"00"		 &"000"&'0'&'0'&'0'&'0'&'1'&'1'&'0'&'1'&"01111"&'1'&'0'&'0'&'1', -- B
		X"00"		 &"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"01111"&'1'&'0'&'0'&'0', -- C
		X"04"		 &"001"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"01111"&'1'&'0'&'0'&'0', -- D
		------------------------------------------------------------------------------
		------------------------------------------------------------------------------
		-- END OF STR INSTRUCTION 
		------------------------------------------------------------------------------
		------------------------------------------------------------------------------
		X"00"		 &"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- E
		X"00"		 &"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- F	
				-- 4
		--NA        MS    MC  IL  PI  PL  TD  TA  TB  MB  FS      MD  RW  MM  MW	
		------------------------------------------------------------------------------
		------------------------------------------------------------------------------
		-- UNCONDITIONAL JMP INSTRUCTION  -  ADDRESS 0x40 -> 0x42
		------------------------------------------------------------------------------
		------------------------------------------------------------------------------
		X"40"		 &"000"&'0'&'0'&'0'&'1'&'0'&'0'&'0'&'0'&"11111"&'1'&'0'&'1'&'0', -- 0
		X"41"		 &"000"&'0'&'1'&'0'&'0'&'0'&'0'&'0'&'0'&"11111"&'0'&'0'&'1'&'0', -- 1
		X"42"		 &"001"&'1'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"11111"&'0'&'0'&'1'&'0', -- 2
		------------------------------------------------------------------------------
		------------------------------------------------------------------------------
		-- END OF JMP INSTRUCTION  
		------------------------------------------------------------------------------
		------------------------------------------------------------------------------
		
		------------------------------------------------------------------------------
		------------------------------------------------------------------------------
		-- BCS INSTRUCTION  -  ADDRESS 0x43 -> 0x47  
		------------------------------------------------------------------------------
		------------------------------------------------------------------------------
		X"4F"		 &"110"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"11111"&'0'&'0'&'1'&'0', -- 3
		X"44"		 &"000"&'0'&'0'&'0'&'1'&'0'&'0'&'0'&'0'&"11111"&'0'&'0'&'1'&'0', -- 4
		X"45"		 &"000"&'0'&'1'&'0'&'0'&'0'&'0'&'0'&'0'&"11111"&'0'&'0'&'1'&'0', -- 5
		X"46"		 &"001"&'1'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"11111"&'0'&'0'&'1'&'0', -- 6
		------------------------------------------------------------------------------
		------------------------------------------------------------------------------
		-- END OF BCS INSTRUCTION 
		------------------------------------------------------------------------------
		------------------------------------------------------------------------------
		------------------------------------------------------------------------------
		
		------------------------------------------------------------------------------
		-- BCC INSTRUCTION  -  ADDRESS 0x48 -> 0x4C  
		------------------------------------------------------------------------------
		------------------------------------------------------------------------------
		X"4F"		 &"010"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"11111"&'0'&'0'&'1'&'0', -- 7
		X"48"		 &"000"&'0'&'0'&'0'&'1'&'0'&'0'&'0'&'0'&"11111"&'0'&'0'&'1'&'0', -- 8
		X"49"		 &"000"&'0'&'1'&'0'&'0'&'0'&'0'&'0'&'0'&"11111"&'0'&'0'&'1'&'0', -- 9
		X"4A"		 &"001"&'1'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"11111"&'0'&'0'&'1'&'0', -- A
		------------------------------------------------------------------------------
		------------------------------------------------------------------------------
		-- END OF BCS INSTRUCTION 
		------------------------------------------------------------------------------
		------------------------------------------------------------------------------
		X"4B"		 &"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"11111"&'0'&'0'&'1'&'0', -- B
		X"4C"		 &"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"11111"&'0'&'0'&'0'&'0', -- C

		X"4D"		 &"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"11111"&'0'&'0'&'0'&'0', -- D
		X"4E"		 &"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"11111"&'0'&'0'&'0'&'0', -- E
		X"4F"		 &"001"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"11111"&'0'&'0'&'0'&'0', -- F
		
				-- 5
		--NA        MS    MC  IL  PI  PL  TD  TA  TB  MB  FS      MD  RW  MM  MW
		x"50"		 &"001"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'1'&"11111"&'1'&'0'&'0'&'0', -- 0
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 1
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 2
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 3
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 4
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 5
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 6
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 7
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 8
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 9
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- A
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- B
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- C
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- D
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- E
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- F
		
				-- 6
		--NA        MS    MC  IL  PI  PL  TD  TA  TB  MB  FS      MD  RW  MM  MW

		X"00" 	 &"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 0		
		X"00"		 &"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 1
		X"00"		 &"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 2
		X"04"		 &"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 3 

		X"64"		 &"001"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"10001"&'0'&'0'&'0'&'0', -- 4
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 5
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 6
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 7
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 8
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 9
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- A
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- B
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- C
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- D
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- E
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- F
		
				-- 7
		--NA        MS    MC  IL  PI  PL  TD  TA  TB  MB  FS      MD  RW  MM  MW
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 0
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 1
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 2
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 3
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 4
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 5
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 6
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 7
		
		x"78" 	 &"001"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'1'&"11111"&'1'&'0'&'1'&'0', -- 8
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 9
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- A
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- B
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- C
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- D
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- E
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- F
		
				-- 8
		--NA        MS    MC  IL  PI  PL  TD  TA  TB  MB  FS      MD  RW  MM  MW
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 0
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 1
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 2
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 3
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 4
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 5
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 6
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 7
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 8
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 9
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- A
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- B
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- C
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- D
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- E
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- F
		
			   -- 9
		--NA        MS    MC  IL  PI  PL  TD  TA  TB  MB  FS      MD  RW  MM  MW
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 0
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 1
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 2
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 3
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 4
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 5
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 6
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 7
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 8
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 9
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- A
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- B
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- C
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- D
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- E
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- F
		
		------------------------------------------------------------------------------
		-- A		DEAL WITH A CURRENT ADD INSTRUCTION
		------------------------------------------------------------------------------		
		--NA        MS    MC  IL  PI  PL  TD  TA  TB  MB  FS      MD  RW  MM  MW
		x"A1"     &"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 0
		x"A2"     &"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 1
		x"FF"		 &"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 2
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 3
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 4
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 5
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 6
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 7
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 8
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 9
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- A
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- B
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- C
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- D
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- E
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- F
		
				-- B
		--NA        MS    MC  IL  PI  PL  TD  TA  TB  MB  FS      MD  RW  MM  MW
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 0
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 1
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 2
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 3
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 4
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 5
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 6
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 7
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 8
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 9
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- A
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- B
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- C
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- D
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- E
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- F
		
				-- C
		--NA        MS    MC  IL  PI  PL  TD  TA  TB  MB  FS      MD  RW  MM  MW
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 0
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 1
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 2
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 3
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 4
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 5
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 6
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 7
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 8
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 9
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- A
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- B
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- C
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- D
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- E
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- F
		
			   -- D
		--NA        MS    MC  IL  PI  PL  TD  TA  TB  MB  FS      MD  RW  MM  MW
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 0
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 1
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 2
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 3
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 4
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 5
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 6
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 7
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 8
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 9
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- A
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- B
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- C
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- D
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- E
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- F
		
			   -- E
		--NA        MS    MC  IL  PI  PL  TD  TA  TB  MB  FS      MD  RW  MM  MW
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 0
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 1
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 2
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 3
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 4
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 5
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 6
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 7
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 8
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 9
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- A
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- B
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- C
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- D
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- E
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- F
		
				-- F
		--NA        MS    MC  IL  PI  PL  TD  TA  TB  MB  FS      MD  RW  MM  MW
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 0
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 1
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 2
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 3
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 4
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 5
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 6
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 7
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 8
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- 9
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- A
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- B
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- C
		"00000000"&"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- D
		x"00"		 &"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0', -- E
		x"ff"     &"000"&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&"00000"&'0'&'0'&'0'&'0' -- F
		);
		
		variable addr : integer;
		variable control_out : std_logic_vector(27 downto 0);
		begin
			addr := conv_integer(IN_CAR);
			control_out := control_mem(addr);
			MW <= control_out(0);
			MM <= control_out(1);
			RW <= control_out(2);
			MD <= control_out(3);
			FUNC_SEL <= control_out(8 downto 4);
			MB <= control_out(9);
			TB <= control_out(10);
			TA <= control_out(11);
			TD <= control_out(12);
			PL <= control_out(13);
			PI <= control_out(14);
			IL <= control_out(15);
			MC <= control_out(16);
			MS_SEL <= control_out(19 downto 17);
			NA <= control_out(27 downto 20);
	end process;
end Behavioral;
